entity VHDL1 is
end entity;

architecture simulation of VHDL1 is
begin

	process is
	begin
	
		report "Hello World";
		wait;
	end process;

end architecture;